module top(output red, output green, output blue);
    assign red   = 0;
    assign green = 1;
    assign blue  = 1;
endmodule